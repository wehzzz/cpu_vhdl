LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY RegAff IS
  PORT (
    Clk : IN STD_LOGIC;
    Reset : IN STD_LOGIC;
    En : IN STD_LOGIC;
    D : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    Q : OUT STD_LOGIC_VECTOR(23 DOWNTO 0)
  );
END ENTITY RegAff;

ARCHITECTURE rtl OF RegAff IS
BEGIN
  PROCESS (Clk, Reset)
  BEGIN
    IF Reset = '1' THEN
      Q <= (OTHERS => '0');
    ELSIF rising_edge(Clk) THEN
      IF En = '1' THEN
        Q <= D(23 DOWNTO 0);
      END IF;
    END IF;
  END PROCESS;
END ARCHITECTURE rtl;